// SISTEMA.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module SISTEMA (
		input  wire        clk_clk,                     //                    clk.clk
		output wire        clk_sdram_clk,               //              clk_sdram.clk
		output wire        ldr_external_interface_sclk, // ldr_external_interface.sclk
		output wire        ldr_external_interface_cs_n, //                       .cs_n
		input  wire        ldr_external_interface_dout, //                       .dout
		output wire        ldr_external_interface_din,  //                       .din
		output wire        pll_locked_export,           //             pll_locked.export
		input  wire        reset_reset_n,               //                  reset.reset_n
		output wire [12:0] sdram_wire_addr,             //             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,               //                       .ba
		output wire        sdram_wire_cas_n,            //                       .cas_n
		output wire        sdram_wire_cke,              //                       .cke
		output wire        sdram_wire_cs_n,             //                       .cs_n
		inout  wire [15:0] sdram_wire_dq,               //                       .dq
		output wire [1:0]  sdram_wire_dqm,              //                       .dqm
		output wire        sdram_wire_ras_n,            //                       .ras_n
		output wire        sdram_wire_we_n              //                       .we_n
	);

	wire          pll_outclk0_clk;                                           // PLL:outclk_0 -> [JTAG_UART:clk, LDR:clock, Procesador1:clk, Procesador2:clk, SDRAM:clk, SRAM1:clk, SRAM2:clk, TIMER:clk, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:PLL_outclk0_clk, rst_controller:clk]
	wire   [31:0] procesador1_data_master_readdata;                          // mm_interconnect_0:Procesador1_data_master_readdata -> Procesador1:d_readdata
	wire          procesador1_data_master_waitrequest;                       // mm_interconnect_0:Procesador1_data_master_waitrequest -> Procesador1:d_waitrequest
	wire          procesador1_data_master_debugaccess;                       // Procesador1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Procesador1_data_master_debugaccess
	wire   [26:0] procesador1_data_master_address;                           // Procesador1:d_address -> mm_interconnect_0:Procesador1_data_master_address
	wire    [3:0] procesador1_data_master_byteenable;                        // Procesador1:d_byteenable -> mm_interconnect_0:Procesador1_data_master_byteenable
	wire          procesador1_data_master_read;                              // Procesador1:d_read -> mm_interconnect_0:Procesador1_data_master_read
	wire          procesador1_data_master_write;                             // Procesador1:d_write -> mm_interconnect_0:Procesador1_data_master_write
	wire   [31:0] procesador1_data_master_writedata;                         // Procesador1:d_writedata -> mm_interconnect_0:Procesador1_data_master_writedata
	wire   [31:0] procesador1_instruction_master_readdata;                   // mm_interconnect_0:Procesador1_instruction_master_readdata -> Procesador1:i_readdata
	wire          procesador1_instruction_master_waitrequest;                // mm_interconnect_0:Procesador1_instruction_master_waitrequest -> Procesador1:i_waitrequest
	wire   [26:0] procesador1_instruction_master_address;                    // Procesador1:i_address -> mm_interconnect_0:Procesador1_instruction_master_address
	wire          procesador1_instruction_master_read;                       // Procesador1:i_read -> mm_interconnect_0:Procesador1_instruction_master_read
	wire   [31:0] procesador2_data_master_readdata;                          // mm_interconnect_0:Procesador2_data_master_readdata -> Procesador2:d_readdata
	wire          procesador2_data_master_waitrequest;                       // mm_interconnect_0:Procesador2_data_master_waitrequest -> Procesador2:d_waitrequest
	wire          procesador2_data_master_debugaccess;                       // Procesador2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Procesador2_data_master_debugaccess
	wire   [26:0] procesador2_data_master_address;                           // Procesador2:d_address -> mm_interconnect_0:Procesador2_data_master_address
	wire    [3:0] procesador2_data_master_byteenable;                        // Procesador2:d_byteenable -> mm_interconnect_0:Procesador2_data_master_byteenable
	wire          procesador2_data_master_read;                              // Procesador2:d_read -> mm_interconnect_0:Procesador2_data_master_read
	wire          procesador2_data_master_write;                             // Procesador2:d_write -> mm_interconnect_0:Procesador2_data_master_write
	wire   [31:0] procesador2_data_master_writedata;                         // Procesador2:d_writedata -> mm_interconnect_0:Procesador2_data_master_writedata
	wire   [31:0] procesador2_instruction_master_readdata;                   // mm_interconnect_0:Procesador2_instruction_master_readdata -> Procesador2:i_readdata
	wire          procesador2_instruction_master_waitrequest;                // mm_interconnect_0:Procesador2_instruction_master_waitrequest -> Procesador2:i_waitrequest
	wire   [26:0] procesador2_instruction_master_address;                    // Procesador2:i_address -> mm_interconnect_0:Procesador2_instruction_master_address
	wire          procesador2_instruction_master_read;                       // Procesador2:i_read -> mm_interconnect_0:Procesador2_instruction_master_read
	wire   [31:0] mm_interconnect_0_ldr_adc_slave_readdata;                  // LDR:readdata -> mm_interconnect_0:LDR_adc_slave_readdata
	wire          mm_interconnect_0_ldr_adc_slave_waitrequest;               // LDR:waitrequest -> mm_interconnect_0:LDR_adc_slave_waitrequest
	wire    [2:0] mm_interconnect_0_ldr_adc_slave_address;                   // mm_interconnect_0:LDR_adc_slave_address -> LDR:address
	wire          mm_interconnect_0_ldr_adc_slave_read;                      // mm_interconnect_0:LDR_adc_slave_read -> LDR:read
	wire          mm_interconnect_0_ldr_adc_slave_write;                     // mm_interconnect_0:LDR_adc_slave_write -> LDR:write
	wire   [31:0] mm_interconnect_0_ldr_adc_slave_writedata;                 // mm_interconnect_0:LDR_adc_slave_writedata -> LDR:writedata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire   [31:0] mm_interconnect_0_procesador1_debug_mem_slave_readdata;    // Procesador1:debug_mem_slave_readdata -> mm_interconnect_0:Procesador1_debug_mem_slave_readdata
	wire          mm_interconnect_0_procesador1_debug_mem_slave_waitrequest; // Procesador1:debug_mem_slave_waitrequest -> mm_interconnect_0:Procesador1_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_procesador1_debug_mem_slave_debugaccess; // mm_interconnect_0:Procesador1_debug_mem_slave_debugaccess -> Procesador1:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_procesador1_debug_mem_slave_address;     // mm_interconnect_0:Procesador1_debug_mem_slave_address -> Procesador1:debug_mem_slave_address
	wire          mm_interconnect_0_procesador1_debug_mem_slave_read;        // mm_interconnect_0:Procesador1_debug_mem_slave_read -> Procesador1:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_procesador1_debug_mem_slave_byteenable;  // mm_interconnect_0:Procesador1_debug_mem_slave_byteenable -> Procesador1:debug_mem_slave_byteenable
	wire          mm_interconnect_0_procesador1_debug_mem_slave_write;       // mm_interconnect_0:Procesador1_debug_mem_slave_write -> Procesador1:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_procesador1_debug_mem_slave_writedata;   // mm_interconnect_0:Procesador1_debug_mem_slave_writedata -> Procesador1:debug_mem_slave_writedata
	wire          mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire   [15:0] mm_interconnect_0_timer_s1_readdata;                       // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire          mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire   [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire          mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire   [15:0] mm_interconnect_0_sdram_s1_readdata;                       // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire          mm_interconnect_0_sdram_s1_waitrequest;                    // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire   [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire          mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire    [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire          mm_interconnect_0_sdram_s1_readdatavalid;                  // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire          mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire   [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire          mm_interconnect_0_sram1_s1_chipselect;                     // mm_interconnect_0:SRAM1_s1_chipselect -> SRAM1:chipselect
	wire  [127:0] mm_interconnect_0_sram1_s1_readdata;                       // SRAM1:readdata -> mm_interconnect_0:SRAM1_s1_readdata
	wire   [12:0] mm_interconnect_0_sram1_s1_address;                        // mm_interconnect_0:SRAM1_s1_address -> SRAM1:address
	wire   [15:0] mm_interconnect_0_sram1_s1_byteenable;                     // mm_interconnect_0:SRAM1_s1_byteenable -> SRAM1:byteenable
	wire          mm_interconnect_0_sram1_s1_write;                          // mm_interconnect_0:SRAM1_s1_write -> SRAM1:write
	wire  [127:0] mm_interconnect_0_sram1_s1_writedata;                      // mm_interconnect_0:SRAM1_s1_writedata -> SRAM1:writedata
	wire          mm_interconnect_0_sram1_s1_clken;                          // mm_interconnect_0:SRAM1_s1_clken -> SRAM1:clken
	wire   [31:0] mm_interconnect_0_procesador2_debug_mem_slave_readdata;    // Procesador2:debug_mem_slave_readdata -> mm_interconnect_0:Procesador2_debug_mem_slave_readdata
	wire          mm_interconnect_0_procesador2_debug_mem_slave_waitrequest; // Procesador2:debug_mem_slave_waitrequest -> mm_interconnect_0:Procesador2_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_procesador2_debug_mem_slave_debugaccess; // mm_interconnect_0:Procesador2_debug_mem_slave_debugaccess -> Procesador2:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_procesador2_debug_mem_slave_address;     // mm_interconnect_0:Procesador2_debug_mem_slave_address -> Procesador2:debug_mem_slave_address
	wire          mm_interconnect_0_procesador2_debug_mem_slave_read;        // mm_interconnect_0:Procesador2_debug_mem_slave_read -> Procesador2:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_procesador2_debug_mem_slave_byteenable;  // mm_interconnect_0:Procesador2_debug_mem_slave_byteenable -> Procesador2:debug_mem_slave_byteenable
	wire          mm_interconnect_0_procesador2_debug_mem_slave_write;       // mm_interconnect_0:Procesador2_debug_mem_slave_write -> Procesador2:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_procesador2_debug_mem_slave_writedata;   // mm_interconnect_0:Procesador2_debug_mem_slave_writedata -> Procesador2:debug_mem_slave_writedata
	wire          mm_interconnect_0_sram2_s1_chipselect;                     // mm_interconnect_0:SRAM2_s1_chipselect -> SRAM2:chipselect
	wire  [127:0] mm_interconnect_0_sram2_s1_readdata;                       // SRAM2:readdata -> mm_interconnect_0:SRAM2_s1_readdata
	wire   [12:0] mm_interconnect_0_sram2_s1_address;                        // mm_interconnect_0:SRAM2_s1_address -> SRAM2:address
	wire   [15:0] mm_interconnect_0_sram2_s1_byteenable;                     // mm_interconnect_0:SRAM2_s1_byteenable -> SRAM2:byteenable
	wire          mm_interconnect_0_sram2_s1_write;                          // mm_interconnect_0:SRAM2_s1_write -> SRAM2:write
	wire  [127:0] mm_interconnect_0_sram2_s1_writedata;                      // mm_interconnect_0:SRAM2_s1_writedata -> SRAM2:writedata
	wire          mm_interconnect_0_sram2_s1_clken;                          // mm_interconnect_0:SRAM2_s1_clken -> SRAM2:clken
	wire   [31:0] procesador1_irq_irq;                                       // irq_mapper:sender_irq -> Procesador1:irq
	wire   [31:0] procesador2_irq_irq;                                       // irq_mapper_001:sender_irq -> Procesador2:irq
	wire          irq_mapper_receiver1_irq;                                  // JTAG_UART:av_irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire          irq_mapper_receiver0_irq;                                  // TIMER:irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [JTAG_UART:rst_n, LDR:reset, Procesador1:reset_n, Procesador2:reset_n, SDRAM:reset_n, SRAM1:reset, SRAM2:reset, TIMER:reset_n, irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:Procesador1_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [Procesador1:reset_req, Procesador2:reset_req, SRAM1:reset_req, SRAM2:reset_req, rst_translator:reset_req_in]
	wire          procesador1_debug_reset_request_reset;                     // Procesador1:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire          procesador2_debug_reset_request_reset;                     // Procesador2:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> PLL:rst

	SISTEMA_JTAG_UART jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	SISTEMA_LDR #(
		.board          ("DE1-SoC"),
		.board_rev      ("Autodetect"),
		.tsclk          (8),
		.numch          (3),
		.max10pllmultby (1),
		.max10plldivby  (1)
	) ldr (
		.clock       (pll_outclk0_clk),                             //                clk.clk
		.reset       (rst_controller_reset_out_reset),              //              reset.reset
		.write       (mm_interconnect_0_ldr_adc_slave_write),       //          adc_slave.write
		.readdata    (mm_interconnect_0_ldr_adc_slave_readdata),    //                   .readdata
		.writedata   (mm_interconnect_0_ldr_adc_slave_writedata),   //                   .writedata
		.address     (mm_interconnect_0_ldr_adc_slave_address),     //                   .address
		.waitrequest (mm_interconnect_0_ldr_adc_slave_waitrequest), //                   .waitrequest
		.read        (mm_interconnect_0_ldr_adc_slave_read),        //                   .read
		.adc_sclk    (ldr_external_interface_sclk),                 // external_interface.export
		.adc_cs_n    (ldr_external_interface_cs_n),                 //                   .export
		.adc_dout    (ldr_external_interface_dout),                 //                   .export
		.adc_din     (ldr_external_interface_din)                   //                   .export
	);

	SISTEMA_PLL pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (pll_outclk0_clk),                    // outclk0.clk
		.outclk_1 (clk_sdram_clk),                      // outclk1.clk
		.locked   (pll_locked_export)                   //  locked.export
	);

	SISTEMA_Procesador1 procesador1 (
		.clk                                 (pll_outclk0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (procesador1_data_master_address),                           //               data_master.address
		.d_byteenable                        (procesador1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (procesador1_data_master_read),                              //                          .read
		.d_readdata                          (procesador1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (procesador1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (procesador1_data_master_write),                             //                          .write
		.d_writedata                         (procesador1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (procesador1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (procesador1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (procesador1_instruction_master_read),                       //                          .read
		.i_readdata                          (procesador1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (procesador1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (procesador1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (procesador1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_procesador1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_procesador1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_procesador1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_procesador1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_procesador1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_procesador1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_procesador1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_procesador1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                           // custom_instruction_master.readra
	);

	SISTEMA_Procesador2 procesador2 (
		.clk                                 (pll_outclk0_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (procesador2_data_master_address),                           //               data_master.address
		.d_byteenable                        (procesador2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (procesador2_data_master_read),                              //                          .read
		.d_readdata                          (procesador2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (procesador2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (procesador2_data_master_write),                             //                          .write
		.d_writedata                         (procesador2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (procesador2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (procesador2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (procesador2_instruction_master_read),                       //                          .read
		.i_readdata                          (procesador2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (procesador2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (procesador2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (procesador2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_procesador2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_procesador2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_procesador2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_procesador2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_procesador2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_procesador2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_procesador2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_procesador2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                           // custom_instruction_master.readra
	);

	SISTEMA_SDRAM sdram (
		.clk            (pll_outclk0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	SISTEMA_SRAM1 sram1 (
		.clk        (pll_outclk0_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_sram1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	SISTEMA_SRAM2 sram2 (
		.clk        (pll_outclk0_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_sram2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	SISTEMA_TIMER timer (
		.clk        (pll_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	SISTEMA_mm_interconnect_0 mm_interconnect_0 (
		.PLL_outclk0_clk                               (pll_outclk0_clk),                                           //                             PLL_outclk0.clk
		.Procesador1_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // Procesador1_reset_reset_bridge_in_reset.reset
		.Procesador1_data_master_address               (procesador1_data_master_address),                           //                 Procesador1_data_master.address
		.Procesador1_data_master_waitrequest           (procesador1_data_master_waitrequest),                       //                                        .waitrequest
		.Procesador1_data_master_byteenable            (procesador1_data_master_byteenable),                        //                                        .byteenable
		.Procesador1_data_master_read                  (procesador1_data_master_read),                              //                                        .read
		.Procesador1_data_master_readdata              (procesador1_data_master_readdata),                          //                                        .readdata
		.Procesador1_data_master_write                 (procesador1_data_master_write),                             //                                        .write
		.Procesador1_data_master_writedata             (procesador1_data_master_writedata),                         //                                        .writedata
		.Procesador1_data_master_debugaccess           (procesador1_data_master_debugaccess),                       //                                        .debugaccess
		.Procesador1_instruction_master_address        (procesador1_instruction_master_address),                    //          Procesador1_instruction_master.address
		.Procesador1_instruction_master_waitrequest    (procesador1_instruction_master_waitrequest),                //                                        .waitrequest
		.Procesador1_instruction_master_read           (procesador1_instruction_master_read),                       //                                        .read
		.Procesador1_instruction_master_readdata       (procesador1_instruction_master_readdata),                   //                                        .readdata
		.Procesador2_data_master_address               (procesador2_data_master_address),                           //                 Procesador2_data_master.address
		.Procesador2_data_master_waitrequest           (procesador2_data_master_waitrequest),                       //                                        .waitrequest
		.Procesador2_data_master_byteenable            (procesador2_data_master_byteenable),                        //                                        .byteenable
		.Procesador2_data_master_read                  (procesador2_data_master_read),                              //                                        .read
		.Procesador2_data_master_readdata              (procesador2_data_master_readdata),                          //                                        .readdata
		.Procesador2_data_master_write                 (procesador2_data_master_write),                             //                                        .write
		.Procesador2_data_master_writedata             (procesador2_data_master_writedata),                         //                                        .writedata
		.Procesador2_data_master_debugaccess           (procesador2_data_master_debugaccess),                       //                                        .debugaccess
		.Procesador2_instruction_master_address        (procesador2_instruction_master_address),                    //          Procesador2_instruction_master.address
		.Procesador2_instruction_master_waitrequest    (procesador2_instruction_master_waitrequest),                //                                        .waitrequest
		.Procesador2_instruction_master_read           (procesador2_instruction_master_read),                       //                                        .read
		.Procesador2_instruction_master_readdata       (procesador2_instruction_master_readdata),                   //                                        .readdata
		.JTAG_UART_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //             JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.JTAG_UART_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.JTAG_UART_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.JTAG_UART_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.LDR_adc_slave_address                         (mm_interconnect_0_ldr_adc_slave_address),                   //                           LDR_adc_slave.address
		.LDR_adc_slave_write                           (mm_interconnect_0_ldr_adc_slave_write),                     //                                        .write
		.LDR_adc_slave_read                            (mm_interconnect_0_ldr_adc_slave_read),                      //                                        .read
		.LDR_adc_slave_readdata                        (mm_interconnect_0_ldr_adc_slave_readdata),                  //                                        .readdata
		.LDR_adc_slave_writedata                       (mm_interconnect_0_ldr_adc_slave_writedata),                 //                                        .writedata
		.LDR_adc_slave_waitrequest                     (mm_interconnect_0_ldr_adc_slave_waitrequest),               //                                        .waitrequest
		.Procesador1_debug_mem_slave_address           (mm_interconnect_0_procesador1_debug_mem_slave_address),     //             Procesador1_debug_mem_slave.address
		.Procesador1_debug_mem_slave_write             (mm_interconnect_0_procesador1_debug_mem_slave_write),       //                                        .write
		.Procesador1_debug_mem_slave_read              (mm_interconnect_0_procesador1_debug_mem_slave_read),        //                                        .read
		.Procesador1_debug_mem_slave_readdata          (mm_interconnect_0_procesador1_debug_mem_slave_readdata),    //                                        .readdata
		.Procesador1_debug_mem_slave_writedata         (mm_interconnect_0_procesador1_debug_mem_slave_writedata),   //                                        .writedata
		.Procesador1_debug_mem_slave_byteenable        (mm_interconnect_0_procesador1_debug_mem_slave_byteenable),  //                                        .byteenable
		.Procesador1_debug_mem_slave_waitrequest       (mm_interconnect_0_procesador1_debug_mem_slave_waitrequest), //                                        .waitrequest
		.Procesador1_debug_mem_slave_debugaccess       (mm_interconnect_0_procesador1_debug_mem_slave_debugaccess), //                                        .debugaccess
		.Procesador2_debug_mem_slave_address           (mm_interconnect_0_procesador2_debug_mem_slave_address),     //             Procesador2_debug_mem_slave.address
		.Procesador2_debug_mem_slave_write             (mm_interconnect_0_procesador2_debug_mem_slave_write),       //                                        .write
		.Procesador2_debug_mem_slave_read              (mm_interconnect_0_procesador2_debug_mem_slave_read),        //                                        .read
		.Procesador2_debug_mem_slave_readdata          (mm_interconnect_0_procesador2_debug_mem_slave_readdata),    //                                        .readdata
		.Procesador2_debug_mem_slave_writedata         (mm_interconnect_0_procesador2_debug_mem_slave_writedata),   //                                        .writedata
		.Procesador2_debug_mem_slave_byteenable        (mm_interconnect_0_procesador2_debug_mem_slave_byteenable),  //                                        .byteenable
		.Procesador2_debug_mem_slave_waitrequest       (mm_interconnect_0_procesador2_debug_mem_slave_waitrequest), //                                        .waitrequest
		.Procesador2_debug_mem_slave_debugaccess       (mm_interconnect_0_procesador2_debug_mem_slave_debugaccess), //                                        .debugaccess
		.SDRAM_s1_address                              (mm_interconnect_0_sdram_s1_address),                        //                                SDRAM_s1.address
		.SDRAM_s1_write                                (mm_interconnect_0_sdram_s1_write),                          //                                        .write
		.SDRAM_s1_read                                 (mm_interconnect_0_sdram_s1_read),                           //                                        .read
		.SDRAM_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                       //                                        .readdata
		.SDRAM_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                      //                                        .writedata
		.SDRAM_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                     //                                        .byteenable
		.SDRAM_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                        .readdatavalid
		.SDRAM_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                    //                                        .waitrequest
		.SDRAM_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                     //                                        .chipselect
		.SRAM1_s1_address                              (mm_interconnect_0_sram1_s1_address),                        //                                SRAM1_s1.address
		.SRAM1_s1_write                                (mm_interconnect_0_sram1_s1_write),                          //                                        .write
		.SRAM1_s1_readdata                             (mm_interconnect_0_sram1_s1_readdata),                       //                                        .readdata
		.SRAM1_s1_writedata                            (mm_interconnect_0_sram1_s1_writedata),                      //                                        .writedata
		.SRAM1_s1_byteenable                           (mm_interconnect_0_sram1_s1_byteenable),                     //                                        .byteenable
		.SRAM1_s1_chipselect                           (mm_interconnect_0_sram1_s1_chipselect),                     //                                        .chipselect
		.SRAM1_s1_clken                                (mm_interconnect_0_sram1_s1_clken),                          //                                        .clken
		.SRAM2_s1_address                              (mm_interconnect_0_sram2_s1_address),                        //                                SRAM2_s1.address
		.SRAM2_s1_write                                (mm_interconnect_0_sram2_s1_write),                          //                                        .write
		.SRAM2_s1_readdata                             (mm_interconnect_0_sram2_s1_readdata),                       //                                        .readdata
		.SRAM2_s1_writedata                            (mm_interconnect_0_sram2_s1_writedata),                      //                                        .writedata
		.SRAM2_s1_byteenable                           (mm_interconnect_0_sram2_s1_byteenable),                     //                                        .byteenable
		.SRAM2_s1_chipselect                           (mm_interconnect_0_sram2_s1_chipselect),                     //                                        .chipselect
		.SRAM2_s1_clken                                (mm_interconnect_0_sram2_s1_clken),                          //                                        .clken
		.TIMER_s1_address                              (mm_interconnect_0_timer_s1_address),                        //                                TIMER_s1.address
		.TIMER_s1_write                                (mm_interconnect_0_timer_s1_write),                          //                                        .write
		.TIMER_s1_readdata                             (mm_interconnect_0_timer_s1_readdata),                       //                                        .readdata
		.TIMER_s1_writedata                            (mm_interconnect_0_timer_s1_writedata),                      //                                        .writedata
		.TIMER_s1_chipselect                           (mm_interconnect_0_timer_s1_chipselect)                      //                                        .chipselect
	);

	SISTEMA_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (procesador1_irq_irq)             //    sender.irq
	);

	SISTEMA_irq_mapper irq_mapper_001 (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (procesador2_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                        // reset_in0.reset
		.reset_in1      (procesador1_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (procesador2_debug_reset_request_reset), // reset_in2.reset
		.clk            (pll_outclk0_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),    //          .reset_req
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                        // reset_in0.reset
		.reset_in1      (procesador1_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (procesador2_debug_reset_request_reset), // reset_in2.reset
		.clk            (),                                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                      // (terminated)
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

endmodule
